// This is a module that implements an AND gate
// assign the AND of a and b to out
module and_gate( 
input a, 
input b, 
output out );