//Design an 8-bit adder.
//There are two 8 bit inputs (in1 and in2) and a single carry-in input bit, cin.
//The outputs are an 8 bit value, [7:0] sum, and a single carry-out output bit, cout.
//The module should utilize the inputs (in1 and in2) and the cin bit to obtain the output sum and cout values.
module adder_8(output [7:0] sum,
                      output cout,
                      input [7:0] in1, in2,
                      input cin);