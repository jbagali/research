//Please finish designing the 8 bit multiplier module (multiplier_8) below.
//There are two 8 bit inputs (A and B) and a 16 bit output (product).
//The module should utilize the inputs (A and B) to determine the output product correctly in its implementation.
module multiplier_8(output [15:0] product, input [7:0] A, B);