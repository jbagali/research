// Design a half adder.
// A half adder adds two bits and produces a sum and carry-out.
// assign the xor of a and b to sum
// assign the and of a and b to cout
module half_adder( 
input a, b,
output cout, sum );