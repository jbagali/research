// Design a counter that counts starting from 1 to 12.

module counter(
    input clk,
    input reset,
    output reg [3:0] q
);