module wire_assign( input in, output out );