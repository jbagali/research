// Create a 100-bit binary adder. The adder adds two 100-bit numbers and a carry-in to produce a 100-bit sum and carry out.

// Hint: There are too many full adders to instantiate, but behavioural code works in this case.

module Adder100( 
    input [99:0] a, b,
    input cin,
    output cout,
    output [99:0] sum );

