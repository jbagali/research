Design a 4-bit adder.
The module below includes the inputs and outputs in the definition.
Please finish the module.

module adder(output [3:0] sum, output cout, input [3:0] in1, in2, input cin);