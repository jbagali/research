`timescale 1 ns/10 ps  // time-unit = 1 ns, precision = 10 ps

module Adder100_tb;

    // duration for each bit = 20 * timescale = 20 * 1 ns  = 20ns
    localparam period = 20;

    reg [99:0] a;
    reg [99:0] b;
    reg cin;

    wire cout;
    wire [99:0] sum;


    integer mismatch_count;

    Adder100 UUT (.a(a), .b(b), .cin(cin), .cout(cout), .sum(sum));

    initial begin
        mismatch_count = 0;

        // Tick 0: Inputs = 100'b1001001001100000010001001010111101000000110000100100001001101011000001001101100011111000001010110011, 100'b0001100000110101110010111101100001101010001101101111110011001100011011011001011000010100001000110010, 1'b1, Generated = cout, sum, Reference = 1'b0, 100'b1010101010010110000100001000011110101010111110010011111100110111011100100110111100001100010011100110
        a = 100'b1001001001100000010001001010111101000000110000100100001001101011000001001101100011111000001010110011; b = 100'b0001100000110101110010111101100001101010001101101111110011001100011011011001011000010100001000110010; cin = 1'b1; // Set input values
        #period;
        if (!(cout === 1'b0 && sum === 100'b1010101010010110000100001000011110101010111110010011111100110111011100100110111100001100010011100110)) begin
            $display("Mismatch at index 0: Inputs = [%b, %b, %b], Generated = [%b, %b], Reference = [%b, %b]", 100'b1001001001100000010001001010111101000000110000100100001001101011000001001101100011111000001010110011, 100'b0001100000110101110010111101100001101010001101101111110011001100011011011001011000010100001000110010, 1'b1, cout, sum, 1'b0, 100'b1010101010010110000100001000011110101010111110010011111100110111011100100110111100001100010011100110);
            mismatch_count = mismatch_count + 1;
        end

        else begin
            $display("Test 0 passed!");
        end

        // Tick 1: Inputs = 100'b0000100100000000011110011111000110000000100000110110101111100110100001101001110110010001111110001011, 100'b1011000011110100011011100110100111101011101101101010001010111111011010100011000101101111101111000110, 1'b0, Generated = cout, sum, Reference = 1'b0, 100'b1011100111110100111010000101101101101100001110100000111010100101111100001100111100000001101101010001
        a = 100'b0000100100000000011110011111000110000000100000110110101111100110100001101001110110010001111110001011; b = 100'b1011000011110100011011100110100111101011101101101010001010111111011010100011000101101111101111000110; cin = 1'b0; // Set input values
        #period;
        if (!(cout === 1'b0 && sum === 100'b1011100111110100111010000101101101101100001110100000111010100101111100001100111100000001101101010001)) begin
            $display("Mismatch at index 1: Inputs = [%b, %b, %b], Generated = [%b, %b], Reference = [%b, %b]", 100'b0000100100000000011110011111000110000000100000110110101111100110100001101001110110010001111110001011, 100'b1011000011110100011011100110100111101011101101101010001010111111011010100011000101101111101111000110, 1'b0, cout, sum, 1'b0, 100'b1011100111110100111010000101101101101100001110100000111010100101111100001100111100000001101101010001);
            mismatch_count = mismatch_count + 1;
        end

        else begin
            $display("Test 1 passed!");
        end

        // Tick 2: Inputs = 100'b1111110011110001100110111001001001100011011100010111101111000010011000101110101010001001111010010101, 100'b0101001110010101011111111011111100101101110111101001001110010011101111000100100110010110101100001001, 1'b0, Generated = cout, sum, Reference = 1'b1, 100'b0101000010000111000110110101000110010001010100000000111101010110000111110011010000100000100110011110
        a = 100'b1111110011110001100110111001001001100011011100010111101111000010011000101110101010001001111010010101; b = 100'b0101001110010101011111111011111100101101110111101001001110010011101111000100100110010110101100001001; cin = 1'b0; // Set input values
        #period;
        if (!(cout === 1'b1 && sum === 100'b0101000010000111000110110101000110010001010100000000111101010110000111110011010000100000100110011110)) begin
            $display("Mismatch at index 2: Inputs = [%b, %b, %b], Generated = [%b, %b], Reference = [%b, %b]", 100'b1111110011110001100110111001001001100011011100010111101111000010011000101110101010001001111010010101, 100'b0101001110010101011111111011111100101101110111101001001110010011101111000100100110010110101100001001, 1'b0, cout, sum, 1'b1, 100'b0101000010000111000110110101000110010001010100000000111101010110000111110011010000100000100110011110);
            mismatch_count = mismatch_count + 1;
        end

        else begin
            $display("Test 2 passed!");
        end

        // Tick 3: Inputs = 100'b1100011110111100100110000011010011111001011100111011101101001011011001110111101000000000001111010111, 100'b0100011100010110010100100111011000101001011100101100001001001010111001101111010001110001010001011110, 1'b1, Generated = cout, sum, Reference = 1'b1, 100'b0000111011010010111010101010101100100010111001100111110110010110010011100110111001110001100000110110
        a = 100'b1100011110111100100110000011010011111001011100111011101101001011011001110111101000000000001111010111; b = 100'b0100011100010110010100100111011000101001011100101100001001001010111001101111010001110001010001011110; cin = 1'b1; // Set input values
        #period;
        if (!(cout === 1'b1 && sum === 100'b0000111011010010111010101010101100100010111001100111110110010110010011100110111001110001100000110110)) begin
            $display("Mismatch at index 3: Inputs = [%b, %b, %b], Generated = [%b, %b], Reference = [%b, %b]", 100'b1100011110111100100110000011010011111001011100111011101101001011011001110111101000000000001111010111, 100'b0100011100010110010100100111011000101001011100101100001001001010111001101111010001110001010001011110, 1'b1, cout, sum, 1'b1, 100'b0000111011010010111010101010101100100010111001100111110110010110010011100110111001110001100000110110);
            mismatch_count = mismatch_count + 1;
        end

        else begin
            $display("Test 3 passed!");
        end

        // Tick 4: Inputs = 100'b0001011011011001010100111001001100110010110110001111011110110001001100011000001010111001110000111000, 100'b0101011000000001110110010001010000000000100000110010000100001001000000101010101111000010001011010101, 1'b0, Generated = cout, sum, Reference = 1'b0, 100'b0110110011011011001011001010011100110011010111000001100010111010001101000010111001111011111100001101
        a = 100'b0001011011011001010100111001001100110010110110001111011110110001001100011000001010111001110000111000; b = 100'b0101011000000001110110010001010000000000100000110010000100001001000000101010101111000010001011010101; cin = 1'b0; // Set input values
        #period;
        if (!(cout === 1'b0 && sum === 100'b0110110011011011001011001010011100110011010111000001100010111010001101000010111001111011111100001101)) begin
            $display("Mismatch at index 4: Inputs = [%b, %b, %b], Generated = [%b, %b], Reference = [%b, %b]", 100'b0001011011011001010100111001001100110010110110001111011110110001001100011000001010111001110000111000, 100'b0101011000000001110110010001010000000000100000110010000100001001000000101010101111000010001011010101, 1'b0, cout, sum, 1'b0, 100'b0110110011011011001011001010011100110011010111000001100010111010001101000010111001111011111100001101);
            mismatch_count = mismatch_count + 1;
        end

        else begin
            $display("Test 4 passed!");
        end

        // Tick 5: Inputs = 100'b0100111011100101100100000001111101001011010001001100000111011100000010011100001101011110000111000000, 100'b0110110101001101001111101011001010011001101011001111111011101011010111110101010100110001010101101010, 1'b1, Generated = cout, sum, Reference = 1'b0, 100'b1011110000110010110011101101000111100100111100011100000011000111011010010001100010001111011100101011
        a = 100'b0100111011100101100100000001111101001011010001001100000111011100000010011100001101011110000111000000; b = 100'b0110110101001101001111101011001010011001101011001111111011101011010111110101010100110001010101101010; cin = 1'b1; // Set input values
        #period;
        if (!(cout === 1'b0 && sum === 100'b1011110000110010110011101101000111100100111100011100000011000111011010010001100010001111011100101011)) begin
            $display("Mismatch at index 5: Inputs = [%b, %b, %b], Generated = [%b, %b], Reference = [%b, %b]", 100'b0100111011100101100100000001111101001011010001001100000111011100000010011100001101011110000111000000, 100'b0110110101001101001111101011001010011001101011001111111011101011010111110101010100110001010101101010, 1'b1, cout, sum, 1'b0, 100'b1011110000110010110011101101000111100100111100011100000011000111011010010001100010001111011100101011);
            mismatch_count = mismatch_count + 1;
        end

        else begin
            $display("Test 5 passed!");
        end

        // Tick 6: Inputs = 100'b0000000101101011101010110001111101010111000001110111111111110100100011101111001111100010101110010110, 100'b0111100010001100001000100100100100011000001010000100101100101000010101110010101110011000010101100101, 1'b0, Generated = cout, sum, Reference = 1'b0, 100'b0111100111110111110011010110100001101111001011111100101100011100111001100001111101111011000011111011
        a = 100'b0000000101101011101010110001111101010111000001110111111111110100100011101111001111100010101110010110; b = 100'b0111100010001100001000100100100100011000001010000100101100101000010101110010101110011000010101100101; cin = 1'b0; // Set input values
        #period;
        if (!(cout === 1'b0 && sum === 100'b0111100111110111110011010110100001101111001011111100101100011100111001100001111101111011000011111011)) begin
            $display("Mismatch at index 6: Inputs = [%b, %b, %b], Generated = [%b, %b], Reference = [%b, %b]", 100'b0000000101101011101010110001111101010111000001110111111111110100100011101111001111100010101110010110, 100'b0111100010001100001000100100100100011000001010000100101100101000010101110010101110011000010101100101, 1'b0, cout, sum, 1'b0, 100'b0111100111110111110011010110100001101111001011111100101100011100111001100001111101111011000011111011);
            mismatch_count = mismatch_count + 1;
        end

        else begin
            $display("Test 6 passed!");
        end

        // Tick 7: Inputs = 100'b0001111000111100101101000101111011111001001000101001011100110000110001010001000001100010010110011010, 100'b0000111101100010010110011010011011000001111000010000011110011011110001100010010001010000100101000100, 1'b1, Generated = cout, sum, Reference = 1'b0, 100'b0010110110011111000011100000010110111011000000111001111011001100100010110011010010110010111011011111
        a = 100'b0001111000111100101101000101111011111001001000101001011100110000110001010001000001100010010110011010; b = 100'b0000111101100010010110011010011011000001111000010000011110011011110001100010010001010000100101000100; cin = 1'b1; // Set input values
        #period;
        if (!(cout === 1'b0 && sum === 100'b0010110110011111000011100000010110111011000000111001111011001100100010110011010010110010111011011111)) begin
            $display("Mismatch at index 7: Inputs = [%b, %b, %b], Generated = [%b, %b], Reference = [%b, %b]", 100'b0001111000111100101101000101111011111001001000101001011100110000110001010001000001100010010110011010, 100'b0000111101100010010110011010011011000001111000010000011110011011110001100010010001010000100101000100, 1'b1, cout, sum, 1'b0, 100'b0010110110011111000011100000010110111011000000111001111011001100100010110011010010110010111011011111);
            mismatch_count = mismatch_count + 1;
        end

        else begin
            $display("Test 7 passed!");
        end

        if (mismatch_count == 0)
            $display("All tests passed!");
        else
            $display("%0d mismatches out of %0d total tests.", mismatch_count, 8);
        $finish;
    end

endmodule