//Design a 4-bit adder.
//There are two 4 bit inputs (in1 and in2) and a single carry-in input bit, cin.
//The adder should utilize the inputs (in1 and in2) and the cin bit to determine the output sum and cout.
//Please finish the module.

module adder(output [3:0] sum, output cout, input [3:0] in1, in2, input cin);