//Please finish designing the 4 bit multiplier module (multiplier_4) below.
//There are two 4 bit inputs (A and B) and an 8 bit output (product).
//The module should utilize the inputs (A and B) to determine the output product correctly in its implementation.
module multiplier_4(output [7:0] product, input [3:0] A, B);