module mac_unit_8(
    input wire [7:0] multiplier,
    input wire [7:0] multiplicand,
    input wire clk,
    input wire rst,
    output reg [15:0] result
);
