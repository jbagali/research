// This is a module that assigns the output to the input
// assign the output out to the input in
module wire_assign( input in, output out );