Design a Verilog module that computes y = x1 * x2 + x3 * x2, where x1, x2, and x3 are inputs, and returns the value as output y.
The module definition below includes the input and output parameters.
Please finish the implementation of this module.

module arithmetic(output [7:0] y, input [7:0] x1, x2, x3);