Design a 4-bit adder.
The module below includes the inputs and outputs in the definition.
The adder should utilize the two 4 bit inputs (in1 and in2) and the cin bit to determine the output sum (4 bits) and cout bit.
Please finish the module.

module adder(output [3:0] sum, output cout, input [3:0] in1, in2, input cin);